`timescale 1ns/1ns
module vga(n_rst, a, d, n_oe, n_we, n_rdy, color_out, hsync_out, vsync_out);

input n_rst;
input [15:0] a; // external address bus
inout [7:0] d; // external data bus
input n_oe, n_we; // memory control signals
inout n_rdy; // memory ready output
output [3:0] color_out; // color output, 2 bits each channel
output hsync_out, vsync_out; // VGA sync lines

/*
Text RAM address: 0xe000 - 0xefff
Color RAM address: 0xf000 - 0xffff
*/

// Pixel clock is generated by a 25.175 MHz generator on board
// In this model 25 MHz is used.
reg pixel_clk;
always begin
    pixel_clk = 1'b0;
    forever #20 pixel_clk = ~pixel_clk;
end

/*
Overall timings:

ssssssbbbppppppp....ppppf
ssssssbbbppppppp....ppppf
     ....       ....
ssssssbbbppppppp....ppppf
FFFFFFFFFFFFFFFF....FFFFF
FFFFFFFFFFFFFFFF....FFFFF
SSSSSSSSSSSSSSSS....SSSSS
BBBBBBBBBBBBBBBB....BBBBB
BBBBBBBBBBBBBBBB....BBBBB

s - horizontal sync pulse (96)
b - horizontal back porch (48)
f - horizontal front porch (16)
p - pixel area (640x480)
F - verical front porch (10)
S - vertical sync pulse (2)
B - vertical back porch (33)
*/

// see /doc/vga.png for pipeline timings

wire [9:0] vy; // line number (total)
wire [9:0] hx; // column number (total)

// column counter
// always enabled
wire n_h_rst;
wire carry_h01;
wire carry_h12;
counter_74161 cnt_h0(
    .clk(pixel_clk),
    .clr_n(n_h_rst),
    .enp(1'b1),
    .ent(1'b1),
    .load_n(1'b1),
    .P(4'b0),
    .Q(hx[3:0]),
    .rco(carry_h01));
counter_74161 cnt_h1(
    .clk(pixel_clk),
    .clr_n(n_h_rst),
    .enp(1'b1),
    .ent(carry_h01),
    .load_n(1'b1),
    .P(4'b0),
    .Q(hx[7:4]),
    .rco(carry_h12));
wire [3:0] cnt_h2_q;
counter_74161 cnt_h2(
    .clk(pixel_clk),
    .clr_n(n_h_rst),
    .enp(1'b1),
    .ent(carry_h12),
    .load_n(1'b1),
    .P(4'b0),
    .Q(cnt_h2_q));
assign hx[9:8] = cnt_h2_q[1:0];

// row counter
// always enabled
wire n_v_rst;
wire v_cnt_ena = 1'b1;
wire carry_v01;
wire carry_v12;
wire v_clk = n_hsync_out;
counter_74161 cnt_v0(
    .clk(v_clk),
    .clr_n(n_v_rst),
    .enp(v_cnt_ena),
    .ent(1'b1),
    .load_n(1'b1),
    .P(4'b0),
    .Q(vy[3:0]),
    .rco(carry_v01));
counter_74161 cnt_v1(
    .clk(v_clk),
    .clr_n(n_v_rst),
    .enp(v_cnt_ena),
    .ent(carry_v01),
    .load_n(1'b1),
    .P(4'b0),
    .Q(vy[7:4]),
    .rco(carry_v12));
wire [3:0] cnt_v2_q;
counter_74161 cnt_v2(
    .clk(v_clk),
    .clr_n(n_v_rst),
    .enp(v_cnt_ena),
    .ent(carry_v12),
    .load_n(1'b1),
    .P(4'b0),
    .Q(cnt_v2_q));
assign vy[9:8] = cnt_v2_q[1:0];

// char column counter: which char to preload
// reset when total column number is just before the visible area
// incremented on the edge of 8 pixels
wire [6:0] ccol = hx[9:3];

wire [4:0] crow = vy[8:4];

wire [11:0] int_a; // internal address bus to read chars when output is active
assign int_a[6:0] = ccol;
assign int_a[11:7] = crow;

// address bus mux: selects address input to the both RAMs
wire a_sel; // 0 - int, 1 - ext
mux_74157 mux_a0(
    .i0(int_a[3:0]),
    .i1(a[3:0]),
    .s(a_sel),
    .n_e(1'b0),
    .z(char_a[3:0]));
mux_74157 mux_a1(
    .i0(int_a[7:4]),
    .i1(a[7:4]),
    .s(a_sel),
    .n_e(1'b0),
    .z(char_a[7:4]));
mux_74157 mux_a2(
    .i0(int_a[11:8]),
    .i1(a[11:8]),
    .s(a_sel),
    .n_e(1'b0),
    .z(char_a[11:8]));

// text RAM
wire [11:0] char_a;
wire [7:0] text_d;
wire n_text_ram_cs;
wire n_text_ram_oe;
wire n_text_ram_we;
async_ram #(.A_WIDTH(12), .INITIAL_VALUE(2)) text_ram(
    .a(char_a),
    .d(text_d),
    .n_cs(n_text_ram_cs),
    .n_oe(n_text_ram_oe),
    .n_we(n_text_ram_we));

// 3-state buffer directing external data bus to the text RAM
wire n_d_to_text_oe;
buffer_74244 buf_char(
    .o(text_d),
    .i(d),
    .n_oe1(n_d_to_text_oe),
    .n_oe2(n_d_to_text_oe));

// color RAM
wire [7:0] color_d;
wire n_color_ram_cs;
wire n_color_ram_oe;
wire n_color_ram_we;
async_ram #(.A_WIDTH(12), .INITIAL_VALUE(8'ha5)) color_ram(
    .a(char_a),
    .d(color_d),
    .n_cs(n_color_ram_cs),
    .n_oe(n_color_ram_oe),
    .n_we(n_color_ram_we));

// 3-state buffer directing external data bus to the color RAM
wire n_d_to_color_oe;
buffer_74244 buf_color(
    .o(color_d),
    .i(d),
    .n_oe1(n_d_to_color_oe),
    .n_oe2(n_d_to_color_oe));

// character generator ROM
wire [14:0] cgrom_a = {3'b0, text_d, vy[3:0]};
wire [7:0] cgrom_d;
rom_28c256 #(.FILENAME("cg.hex")) cg_rom(
    .a(cgrom_a),
    .d(cgrom_d),
    .n_cs(1'b0),
    .n_oe(1'b0));

// registers to preload 8 pixels of the characters and color
wire buf_clk = ~hx[2];
wire [7:0] stored_pixel;
register_74273 reg_char(
          .q(stored_pixel),
          .d(cgrom_d),
          .n_mr(n_rst),
          .cp(buf_clk));

wire [7:0] stored_color;
register_74273 reg_color(
        .q(stored_color),
        .d(color_d),
        .n_mr(n_rst),
        .cp(buf_clk));

// mux to select a pixel from the preloaded row
wire n_pixel_ena;
wire pixel_out;
mux_74151 mux_pixel(
    .n_g(1'b0),
    .d(stored_pixel),
    .a(hx[0]),
    .b(hx[1]),
    .c(hx[2]),
    .y(pixel_out));

// mux to select bg or fg color based on pixel
mux_74157 mux_color(
    .i0(stored_color[7:4]),
    .i1(stored_color[3:0]),
    .s(pixel_out),
    .n_e(n_pixel_ena),
    .z(color_out));

wire n_hsync_out;

vga_ctrl ctrl(
    .a_sel(a_sel),
    .n_text_ram_cs(n_text_ram_cs),
    .n_text_ram_oe(n_text_ram_oe),
    .n_text_ram_we(n_text_ram_we),
    .n_d_to_text_oe(n_d_to_text_oe),
    .n_color_ram_cs(n_color_ram_cs),
    .n_color_ram_oe(n_color_ram_oe),
    .n_color_ram_we(n_color_ram_we),
    .n_d_to_color_oe(n_d_to_color_oe),
    .n_pixel_ena(n_pixel_ena),
    .n_h_rst(n_h_rst),
    .n_v_rst(n_v_rst),
    .n_hsync_out(n_hsync_out),
    .hsync_out(hsync_out),
    .vsync_out(vsync_out),
    .n_rdy(n_rdy),
    .n_rst(n_rst),
    .a(a),
    .n_we(n_we),
    .n_oe(n_oe),
    .vy(vy),
    .hx(hx));

endmodule
